package decisionTree_fixpt_pkg;
  typedef  logic  [12:0] vector_of_unsigned_logic_13;
endpackage: decisionTree_fixpt_pkg
